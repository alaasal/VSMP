module INPUTREG();
endmodule