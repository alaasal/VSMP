module OUTPUTREG();
endmodule